package shared_pkg;
    int period;
    int count;
    bit have_address;
    logic [10:0] curr_op;
endpackage